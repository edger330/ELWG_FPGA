library verilog;
use verilog.vl_types.all;
entity PU4 is
    port(
        sys_clk         : in     vl_logic;
        sys_rst_n       : in     vl_logic;
        mode            : in     vl_logic;
        SUM_select      : in     vl_logic_vector(2 downto 0);
        Y_Init          : in     vl_logic_vector(31 downto 0);
        SUM_valid       : in     vl_logic;
        SUM_start       : in     vl_logic;
        p_mx_0          : in     vl_logic_vector(31 downto 0);
        p_my_0          : in     vl_logic_vector(31 downto 0);
        p_mm_0          : in     vl_logic_vector(31 downto 0);
        p_mx_1          : in     vl_logic_vector(31 downto 0);
        p_my_1          : in     vl_logic_vector(31 downto 0);
        p_mm_1          : in     vl_logic_vector(31 downto 0);
        p_mx_2          : in     vl_logic_vector(31 downto 0);
        p_my_2          : in     vl_logic_vector(31 downto 0);
        p_mm_2          : in     vl_logic_vector(31 downto 0);
        p_mx_3          : in     vl_logic_vector(31 downto 0);
        p_my_3          : in     vl_logic_vector(31 downto 0);
        p_mm_3          : in     vl_logic_vector(31 downto 0);
        lambda1_0       : in     vl_logic_vector(31 downto 0);
        lambda2_0       : in     vl_logic_vector(31 downto 0);
        lambda1_1       : in     vl_logic_vector(31 downto 0);
        lambda2_1       : in     vl_logic_vector(31 downto 0);
        lambda1_2       : in     vl_logic_vector(31 downto 0);
        lambda2_2       : in     vl_logic_vector(31 downto 0);
        lambda1_3       : in     vl_logic_vector(31 downto 0);
        lambda2_3       : in     vl_logic_vector(31 downto 0);
        H_in            : in     vl_logic_vector(7 downto 0);
        R_in_0          : in     vl_logic_vector(7 downto 0);
        R_in_1          : in     vl_logic_vector(7 downto 0);
        R_in_2          : in     vl_logic_vector(7 downto 0);
        R_in_3          : in     vl_logic_vector(7 downto 0);
        Init_in         : in     vl_logic;
        SUM_out         : out    vl_logic_vector(31 downto 0)
    );
end PU4;
