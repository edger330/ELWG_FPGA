library verilog;
use verilog.vl_types.all;
entity save_send is
    generic(
        PE_NUM          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        ADDR_R          : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_H          : vl_logic_vector(0 to 8) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_QIDC       : vl_logic_vector(0 to 8) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        IDLE            : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        GET_PKT_INFO    : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        GET_R           : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        GET_H           : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        GET_QIDC        : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        WAIT_VLD        : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        PREPARE         : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CALCULATE       : vl_logic_vector(0 to 8) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DONE            : vl_logic_vector(0 to 8) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CAL_IDLE        : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        S0              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        S1              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        S2              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        S3              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        S4              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        S5              : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WAIT_6          : vl_logic_vector(0 to 8) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CAL_DONE        : vl_logic_vector(0 to 8) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        sys_clk         : in     vl_logic;
        sys_rst_n       : in     vl_logic;
        matrix_memory_sop: in     vl_logic;
        matrix_memory_eop: in     vl_logic;
        matrix_memory_vld: in     vl_logic;
        matrix_memory_data: in     vl_logic_vector(31 downto 0);
        vld             : in     vl_logic;
        M_write         : in     vl_logic_vector(31 downto 0);
        X_write         : in     vl_logic_vector(31 downto 0);
        init_out        : in     vl_logic;
        pkt_receive_enable: out    vl_logic;
        ram_out         : out    vl_logic_vector(31 downto 0);
        q               : out    vl_logic_vector(7 downto 0);
        i               : out    vl_logic_vector(7 downto 0);
        r               : out    vl_logic_vector(7 downto 0);
        h               : out    vl_logic_vector(7 downto 0);
        M_read          : out    vl_logic_vector(31 downto 0);
        X_read          : out    vl_logic_vector(31 downto 0);
        parameter_vld   : out    vl_logic;
        en_sum          : out    vl_logic;
        mode            : out    vl_logic;
        sum_select      : out    vl_logic_vector(5 downto 0);
        sum_vld         : out    vl_logic;
        y_initial       : out    vl_logic_vector(31 downto 0);
        init            : out    vl_logic;
        head            : out    vl_logic_vector(63 downto 0);
        pe_cnt          : out    vl_logic_vector(5 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PE_NUM : constant is 1;
    attribute mti_svvh_generic_type of ADDR_R : constant is 1;
    attribute mti_svvh_generic_type of ADDR_H : constant is 1;
    attribute mti_svvh_generic_type of ADDR_QIDC : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of GET_PKT_INFO : constant is 1;
    attribute mti_svvh_generic_type of GET_R : constant is 1;
    attribute mti_svvh_generic_type of GET_H : constant is 1;
    attribute mti_svvh_generic_type of GET_QIDC : constant is 1;
    attribute mti_svvh_generic_type of WAIT_VLD : constant is 1;
    attribute mti_svvh_generic_type of PREPARE : constant is 1;
    attribute mti_svvh_generic_type of CALCULATE : constant is 1;
    attribute mti_svvh_generic_type of DONE : constant is 1;
    attribute mti_svvh_generic_type of CAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of S0 : constant is 1;
    attribute mti_svvh_generic_type of S1 : constant is 1;
    attribute mti_svvh_generic_type of S2 : constant is 1;
    attribute mti_svvh_generic_type of S3 : constant is 1;
    attribute mti_svvh_generic_type of S4 : constant is 1;
    attribute mti_svvh_generic_type of S5 : constant is 1;
    attribute mti_svvh_generic_type of WAIT_6 : constant is 1;
    attribute mti_svvh_generic_type of CAL_DONE : constant is 1;
end save_send;
