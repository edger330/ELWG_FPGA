library verilog;
use verilog.vl_types.all;
entity matrix_memory is
    generic(
        ADDR_HEAD0      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_HEAD1      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        ADDR_HEAD2      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        ADDR_HEAD3      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        ADDR_HEAD4      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        ADDR_HEAD5      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        ADDR_Y_INITIAL  : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        ADDR_LEN        : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        ADDR_HAP_ID     : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        ADDR_P0         : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        ADDR_P1         : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        ADDR_P2         : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ADDR_P3         : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1);
        ADDR_P4         : vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        ADDR_P5         : vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        ADDR_P6         : vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ADDR_RH         : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        ADDR_M_R0       : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_X_R0       : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        ADDR_Y_R0       : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        ADDR_M_R1       : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_X_R1       : vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        ADDR_Y_R1       : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        D               : real    := 0.200000
    );
    port(
        matrix_memory_sop: in     vl_logic;
        matrix_memory_eop: in     vl_logic;
        matrix_memory_vld: in     vl_logic;
        matrix_memory_data: in     vl_logic_vector(31 downto 0);
        m_i_j           : in     vl_logic_vector(31 downto 0);
        x_i_j           : in     vl_logic_vector(31 downto 0);
        y_i_j           : in     vl_logic_vector(31 downto 0);
        vld             : in     vl_logic;
        sys_clk         : in     vl_logic;
        sys_rst         : in     vl_logic;
        number          : in     vl_logic_vector(4 downto 0);
        symbol          : out    vl_logic_vector(4 downto 0);
        p_mx            : out    vl_logic_vector(31 downto 0);
        p_my            : out    vl_logic_vector(31 downto 0);
        p_xx_yy         : out    vl_logic_vector(31 downto 0);
        p_xm_ym         : out    vl_logic_vector(31 downto 0);
        p_mm            : out    vl_logic_vector(31 downto 0);
        m_i1_j1         : out    vl_logic_vector(31 downto 0);
        m_i1_j          : out    vl_logic_vector(31 downto 0);
        x_i1_j1         : out    vl_logic_vector(31 downto 0);
        x_i1_j          : out    vl_logic_vector(31 downto 0);
        y_i1_j1         : out    vl_logic_vector(31 downto 0);
        counter_out_ready_ok: out    vl_logic_vector(3 downto 0);
        counter_row_scan1: out    vl_logic_vector(8 downto 0);
        counter_col_scan1: out    vl_logic_vector(6 downto 0);
        read_len_ok     : out    vl_logic_vector(7 downto 0);
        counter_sum     : out    vl_logic_vector(8 downto 0);
        en_counter_sum  : out    vl_logic;
        busy            : out    vl_logic;
        hap_length      : out    vl_logic_vector(15 downto 0);
        head_read_hap_id: out    vl_logic_vector(95 downto 0);
        counter_head    : out    vl_logic_vector(4 downto 0);
        \signal\        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ADDR_HEAD0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEAD1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEAD2 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEAD3 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEAD4 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEAD5 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_Y_INITIAL : constant is 1;
    attribute mti_svvh_generic_type of ADDR_LEN : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HAP_ID : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P2 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P3 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P4 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P5 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_P6 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_RH : constant is 1;
    attribute mti_svvh_generic_type of ADDR_M_R0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_X_R0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_Y_R0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_M_R1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_X_R1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_Y_R1 : constant is 1;
    attribute mti_svvh_generic_type of D : constant is 1;
end matrix_memory;
