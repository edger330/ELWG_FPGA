library verilog;
use verilog.vl_types.all;
entity PU32 is
    port(
        sys_clk         : in     vl_logic;
        sys_rst_n       : in     vl_logic;
        mode            : in     vl_logic;
        SUM_select      : in     vl_logic_vector(4 downto 0);
        Y_Init          : in     vl_logic_vector(31 downto 0);
        SUM_valid       : in     vl_logic;
        SUM_start       : in     vl_logic;
        p_mx_0          : in     vl_logic_vector(31 downto 0);
        p_my_0          : in     vl_logic_vector(31 downto 0);
        p_mm_0          : in     vl_logic_vector(31 downto 0);
        p_mx_1          : in     vl_logic_vector(31 downto 0);
        p_my_1          : in     vl_logic_vector(31 downto 0);
        p_mm_1          : in     vl_logic_vector(31 downto 0);
        p_mx_2          : in     vl_logic_vector(31 downto 0);
        p_my_2          : in     vl_logic_vector(31 downto 0);
        p_mm_2          : in     vl_logic_vector(31 downto 0);
        p_mx_3          : in     vl_logic_vector(31 downto 0);
        p_my_3          : in     vl_logic_vector(31 downto 0);
        p_mm_3          : in     vl_logic_vector(31 downto 0);
        p_mx_4          : in     vl_logic_vector(31 downto 0);
        p_my_4          : in     vl_logic_vector(31 downto 0);
        p_mm_4          : in     vl_logic_vector(31 downto 0);
        p_mx_5          : in     vl_logic_vector(31 downto 0);
        p_my_5          : in     vl_logic_vector(31 downto 0);
        p_mm_5          : in     vl_logic_vector(31 downto 0);
        p_mx_6          : in     vl_logic_vector(31 downto 0);
        p_my_6          : in     vl_logic_vector(31 downto 0);
        p_mm_6          : in     vl_logic_vector(31 downto 0);
        p_mx_7          : in     vl_logic_vector(31 downto 0);
        p_my_7          : in     vl_logic_vector(31 downto 0);
        p_mm_7          : in     vl_logic_vector(31 downto 0);
        p_mx_8          : in     vl_logic_vector(31 downto 0);
        p_my_8          : in     vl_logic_vector(31 downto 0);
        p_mm_8          : in     vl_logic_vector(31 downto 0);
        p_mx_9          : in     vl_logic_vector(31 downto 0);
        p_my_9          : in     vl_logic_vector(31 downto 0);
        p_mm_9          : in     vl_logic_vector(31 downto 0);
        p_mx_10         : in     vl_logic_vector(31 downto 0);
        p_my_10         : in     vl_logic_vector(31 downto 0);
        p_mm_10         : in     vl_logic_vector(31 downto 0);
        p_mx_11         : in     vl_logic_vector(31 downto 0);
        p_my_11         : in     vl_logic_vector(31 downto 0);
        p_mm_11         : in     vl_logic_vector(31 downto 0);
        p_mx_12         : in     vl_logic_vector(31 downto 0);
        p_my_12         : in     vl_logic_vector(31 downto 0);
        p_mm_12         : in     vl_logic_vector(31 downto 0);
        p_mx_13         : in     vl_logic_vector(31 downto 0);
        p_my_13         : in     vl_logic_vector(31 downto 0);
        p_mm_13         : in     vl_logic_vector(31 downto 0);
        p_mx_14         : in     vl_logic_vector(31 downto 0);
        p_my_14         : in     vl_logic_vector(31 downto 0);
        p_mm_14         : in     vl_logic_vector(31 downto 0);
        p_mx_15         : in     vl_logic_vector(31 downto 0);
        p_my_15         : in     vl_logic_vector(31 downto 0);
        p_mm_15         : in     vl_logic_vector(31 downto 0);
        p_mx_16         : in     vl_logic_vector(31 downto 0);
        p_my_16         : in     vl_logic_vector(31 downto 0);
        p_mm_16         : in     vl_logic_vector(31 downto 0);
        p_mx_17         : in     vl_logic_vector(31 downto 0);
        p_my_17         : in     vl_logic_vector(31 downto 0);
        p_mm_17         : in     vl_logic_vector(31 downto 0);
        p_mx_18         : in     vl_logic_vector(31 downto 0);
        p_my_18         : in     vl_logic_vector(31 downto 0);
        p_mm_18         : in     vl_logic_vector(31 downto 0);
        p_mx_19         : in     vl_logic_vector(31 downto 0);
        p_my_19         : in     vl_logic_vector(31 downto 0);
        p_mm_19         : in     vl_logic_vector(31 downto 0);
        p_mx_20         : in     vl_logic_vector(31 downto 0);
        p_my_20         : in     vl_logic_vector(31 downto 0);
        p_mm_20         : in     vl_logic_vector(31 downto 0);
        p_mx_21         : in     vl_logic_vector(31 downto 0);
        p_my_21         : in     vl_logic_vector(31 downto 0);
        p_mm_21         : in     vl_logic_vector(31 downto 0);
        p_mx_22         : in     vl_logic_vector(31 downto 0);
        p_my_22         : in     vl_logic_vector(31 downto 0);
        p_mm_22         : in     vl_logic_vector(31 downto 0);
        p_mx_23         : in     vl_logic_vector(31 downto 0);
        p_my_23         : in     vl_logic_vector(31 downto 0);
        p_mm_23         : in     vl_logic_vector(31 downto 0);
        p_mx_24         : in     vl_logic_vector(31 downto 0);
        p_my_24         : in     vl_logic_vector(31 downto 0);
        p_mm_24         : in     vl_logic_vector(31 downto 0);
        p_mx_25         : in     vl_logic_vector(31 downto 0);
        p_my_25         : in     vl_logic_vector(31 downto 0);
        p_mm_25         : in     vl_logic_vector(31 downto 0);
        p_mx_26         : in     vl_logic_vector(31 downto 0);
        p_my_26         : in     vl_logic_vector(31 downto 0);
        p_mm_26         : in     vl_logic_vector(31 downto 0);
        p_mx_27         : in     vl_logic_vector(31 downto 0);
        p_my_27         : in     vl_logic_vector(31 downto 0);
        p_mm_27         : in     vl_logic_vector(31 downto 0);
        p_mx_28         : in     vl_logic_vector(31 downto 0);
        p_my_28         : in     vl_logic_vector(31 downto 0);
        p_mm_28         : in     vl_logic_vector(31 downto 0);
        p_mx_29         : in     vl_logic_vector(31 downto 0);
        p_my_29         : in     vl_logic_vector(31 downto 0);
        p_mm_29         : in     vl_logic_vector(31 downto 0);
        p_mx_30         : in     vl_logic_vector(31 downto 0);
        p_my_30         : in     vl_logic_vector(31 downto 0);
        p_mm_30         : in     vl_logic_vector(31 downto 0);
        p_mx_31         : in     vl_logic_vector(31 downto 0);
        p_my_31         : in     vl_logic_vector(31 downto 0);
        p_mm_31         : in     vl_logic_vector(31 downto 0);
        lambda1_0       : in     vl_logic_vector(31 downto 0);
        lambda2_0       : in     vl_logic_vector(31 downto 0);
        lambda1_1       : in     vl_logic_vector(31 downto 0);
        lambda2_1       : in     vl_logic_vector(31 downto 0);
        lambda1_2       : in     vl_logic_vector(31 downto 0);
        lambda2_2       : in     vl_logic_vector(31 downto 0);
        lambda1_3       : in     vl_logic_vector(31 downto 0);
        lambda2_3       : in     vl_logic_vector(31 downto 0);
        lambda1_4       : in     vl_logic_vector(31 downto 0);
        lambda2_4       : in     vl_logic_vector(31 downto 0);
        lambda1_5       : in     vl_logic_vector(31 downto 0);
        lambda2_5       : in     vl_logic_vector(31 downto 0);
        lambda1_6       : in     vl_logic_vector(31 downto 0);
        lambda2_6       : in     vl_logic_vector(31 downto 0);
        lambda1_7       : in     vl_logic_vector(31 downto 0);
        lambda2_7       : in     vl_logic_vector(31 downto 0);
        lambda1_8       : in     vl_logic_vector(31 downto 0);
        lambda2_8       : in     vl_logic_vector(31 downto 0);
        lambda1_9       : in     vl_logic_vector(31 downto 0);
        lambda2_9       : in     vl_logic_vector(31 downto 0);
        lambda1_10      : in     vl_logic_vector(31 downto 0);
        lambda2_10      : in     vl_logic_vector(31 downto 0);
        lambda1_11      : in     vl_logic_vector(31 downto 0);
        lambda2_11      : in     vl_logic_vector(31 downto 0);
        lambda1_12      : in     vl_logic_vector(31 downto 0);
        lambda2_12      : in     vl_logic_vector(31 downto 0);
        lambda1_13      : in     vl_logic_vector(31 downto 0);
        lambda2_13      : in     vl_logic_vector(31 downto 0);
        lambda1_14      : in     vl_logic_vector(31 downto 0);
        lambda2_14      : in     vl_logic_vector(31 downto 0);
        lambda1_15      : in     vl_logic_vector(31 downto 0);
        lambda2_15      : in     vl_logic_vector(31 downto 0);
        lambda1_16      : in     vl_logic_vector(31 downto 0);
        lambda2_16      : in     vl_logic_vector(31 downto 0);
        lambda1_17      : in     vl_logic_vector(31 downto 0);
        lambda2_17      : in     vl_logic_vector(31 downto 0);
        lambda1_18      : in     vl_logic_vector(31 downto 0);
        lambda2_18      : in     vl_logic_vector(31 downto 0);
        lambda1_19      : in     vl_logic_vector(31 downto 0);
        lambda2_19      : in     vl_logic_vector(31 downto 0);
        lambda1_20      : in     vl_logic_vector(31 downto 0);
        lambda2_20      : in     vl_logic_vector(31 downto 0);
        lambda1_21      : in     vl_logic_vector(31 downto 0);
        lambda2_21      : in     vl_logic_vector(31 downto 0);
        lambda1_22      : in     vl_logic_vector(31 downto 0);
        lambda2_22      : in     vl_logic_vector(31 downto 0);
        lambda1_23      : in     vl_logic_vector(31 downto 0);
        lambda2_23      : in     vl_logic_vector(31 downto 0);
        lambda1_24      : in     vl_logic_vector(31 downto 0);
        lambda2_24      : in     vl_logic_vector(31 downto 0);
        lambda1_25      : in     vl_logic_vector(31 downto 0);
        lambda2_25      : in     vl_logic_vector(31 downto 0);
        lambda1_26      : in     vl_logic_vector(31 downto 0);
        lambda2_26      : in     vl_logic_vector(31 downto 0);
        lambda1_27      : in     vl_logic_vector(31 downto 0);
        lambda2_27      : in     vl_logic_vector(31 downto 0);
        lambda1_28      : in     vl_logic_vector(31 downto 0);
        lambda2_28      : in     vl_logic_vector(31 downto 0);
        lambda1_29      : in     vl_logic_vector(31 downto 0);
        lambda2_29      : in     vl_logic_vector(31 downto 0);
        lambda1_30      : in     vl_logic_vector(31 downto 0);
        lambda2_30      : in     vl_logic_vector(31 downto 0);
        lambda1_31      : in     vl_logic_vector(31 downto 0);
        lambda2_31      : in     vl_logic_vector(31 downto 0);
        H_in            : in     vl_logic_vector(7 downto 0);
        R_in_0          : in     vl_logic_vector(7 downto 0);
        R_in_1          : in     vl_logic_vector(7 downto 0);
        R_in_2          : in     vl_logic_vector(7 downto 0);
        R_in_3          : in     vl_logic_vector(7 downto 0);
        R_in_4          : in     vl_logic_vector(7 downto 0);
        R_in_5          : in     vl_logic_vector(7 downto 0);
        R_in_6          : in     vl_logic_vector(7 downto 0);
        R_in_7          : in     vl_logic_vector(7 downto 0);
        R_in_8          : in     vl_logic_vector(7 downto 0);
        R_in_9          : in     vl_logic_vector(7 downto 0);
        R_in_10         : in     vl_logic_vector(7 downto 0);
        R_in_11         : in     vl_logic_vector(7 downto 0);
        R_in_12         : in     vl_logic_vector(7 downto 0);
        R_in_13         : in     vl_logic_vector(7 downto 0);
        R_in_14         : in     vl_logic_vector(7 downto 0);
        R_in_15         : in     vl_logic_vector(7 downto 0);
        R_in_16         : in     vl_logic_vector(7 downto 0);
        R_in_17         : in     vl_logic_vector(7 downto 0);
        R_in_18         : in     vl_logic_vector(7 downto 0);
        R_in_19         : in     vl_logic_vector(7 downto 0);
        R_in_20         : in     vl_logic_vector(7 downto 0);
        R_in_21         : in     vl_logic_vector(7 downto 0);
        R_in_22         : in     vl_logic_vector(7 downto 0);
        R_in_23         : in     vl_logic_vector(7 downto 0);
        R_in_24         : in     vl_logic_vector(7 downto 0);
        R_in_25         : in     vl_logic_vector(7 downto 0);
        R_in_26         : in     vl_logic_vector(7 downto 0);
        R_in_27         : in     vl_logic_vector(7 downto 0);
        R_in_28         : in     vl_logic_vector(7 downto 0);
        R_in_29         : in     vl_logic_vector(7 downto 0);
        R_in_30         : in     vl_logic_vector(7 downto 0);
        R_in_31         : in     vl_logic_vector(7 downto 0);
        Init_in         : in     vl_logic;
        SUM_out         : out    vl_logic_vector(31 downto 0)
    );
end PU32;
